module delay(in,out);
parameter n_delay = 5;//maximum n_delay is 80

input in /*synthesis keep*/;
output out /*synthesis keep*/; 
//synthesis keep = 1;
wire [158:0] internal_wire /*synthesis keep*/;

// four inverters in chain
assign out = ~internal_wire[n_delay*2-2];

assign internal_wire[0] = ~in;
assign internal_wire[1] = ~internal_wire[0];
assign internal_wire[2] = ~internal_wire[1];
assign internal_wire[3] = ~internal_wire[2];
assign internal_wire[4] = ~internal_wire[3];
assign internal_wire[5] = ~internal_wire[4];
assign internal_wire[6] = ~internal_wire[5];
assign internal_wire[7] = ~internal_wire[6];
assign internal_wire[8] = ~internal_wire[7];
assign internal_wire[9] = ~internal_wire[8];
assign internal_wire[10] = ~internal_wire[9];
assign internal_wire[11] = ~internal_wire[10];
assign internal_wire[12] = ~internal_wire[11];
assign internal_wire[13] = ~internal_wire[12];
assign internal_wire[14] = ~internal_wire[13];
assign internal_wire[15] = ~internal_wire[14];
assign internal_wire[16] = ~internal_wire[15];
assign internal_wire[17] = ~internal_wire[16];
assign internal_wire[18] = ~internal_wire[17];
assign internal_wire[19] = ~internal_wire[18];
assign internal_wire[20] = ~internal_wire[19];
assign internal_wire[21] = ~internal_wire[20];
assign internal_wire[22] = ~internal_wire[21];
assign internal_wire[23] = ~internal_wire[22];
assign internal_wire[24] = ~internal_wire[23];
assign internal_wire[25] = ~internal_wire[24];
assign internal_wire[26] = ~internal_wire[25];
assign internal_wire[27] = ~internal_wire[26];
assign internal_wire[28] = ~internal_wire[27];
assign internal_wire[29] = ~internal_wire[28];
assign internal_wire[30] = ~internal_wire[29];
assign internal_wire[31] = ~internal_wire[30];
assign internal_wire[32] = ~internal_wire[31];
assign internal_wire[33] = ~internal_wire[32];
assign internal_wire[34] = ~internal_wire[33];
assign internal_wire[35] = ~internal_wire[34];
assign internal_wire[36] = ~internal_wire[35];
assign internal_wire[37] = ~internal_wire[36];
assign internal_wire[38] = ~internal_wire[37];
assign internal_wire[39] = ~internal_wire[38];
assign internal_wire[40] = ~internal_wire[39];
assign internal_wire[41] = ~internal_wire[40];
assign internal_wire[42] = ~internal_wire[41];
assign internal_wire[43] = ~internal_wire[42];
assign internal_wire[44] = ~internal_wire[43];
assign internal_wire[45] = ~internal_wire[44];
assign internal_wire[46] = ~internal_wire[45];
assign internal_wire[47] = ~internal_wire[46];
assign internal_wire[48] = ~internal_wire[47];
assign internal_wire[49] = ~internal_wire[48];
assign internal_wire[50] = ~internal_wire[49];
assign internal_wire[51] = ~internal_wire[50];
assign internal_wire[52] = ~internal_wire[51];
assign internal_wire[53] = ~internal_wire[52];
assign internal_wire[54] = ~internal_wire[53];
assign internal_wire[55] = ~internal_wire[54];
assign internal_wire[56] = ~internal_wire[55];
assign internal_wire[57] = ~internal_wire[56];
assign internal_wire[58] = ~internal_wire[57];
assign internal_wire[59] = ~internal_wire[58];
assign internal_wire[60] = ~internal_wire[59];
assign internal_wire[61] = ~internal_wire[60];
assign internal_wire[62] = ~internal_wire[61];
assign internal_wire[63] = ~internal_wire[62];
assign internal_wire[64] = ~internal_wire[63];
assign internal_wire[65] = ~internal_wire[64];
assign internal_wire[66] = ~internal_wire[65];
assign internal_wire[67] = ~internal_wire[66];
assign internal_wire[68] = ~internal_wire[67];
assign internal_wire[69] = ~internal_wire[68];
assign internal_wire[70] = ~internal_wire[69];
assign internal_wire[71] = ~internal_wire[70];
assign internal_wire[72] = ~internal_wire[71];
assign internal_wire[73] = ~internal_wire[72];
assign internal_wire[74] = ~internal_wire[73];
assign internal_wire[75] = ~internal_wire[74];
assign internal_wire[76] = ~internal_wire[75];
assign internal_wire[77] = ~internal_wire[76];
assign internal_wire[78] = ~internal_wire[77];
assign internal_wire[79] = ~internal_wire[78];
assign internal_wire[80] = ~internal_wire[79];
assign internal_wire[81] = ~internal_wire[80];
assign internal_wire[82] = ~internal_wire[81];
assign internal_wire[83] = ~internal_wire[82];
assign internal_wire[84] = ~internal_wire[83];
assign internal_wire[85] = ~internal_wire[84];
assign internal_wire[86] = ~internal_wire[85];
assign internal_wire[87] = ~internal_wire[86];
assign internal_wire[88] = ~internal_wire[87];
assign internal_wire[89] = ~internal_wire[88];
assign internal_wire[90] = ~internal_wire[89];
assign internal_wire[91] = ~internal_wire[90];
assign internal_wire[92] = ~internal_wire[91];
assign internal_wire[93] = ~internal_wire[92];
assign internal_wire[94] = ~internal_wire[93];
assign internal_wire[95] = ~internal_wire[94];
assign internal_wire[96] = ~internal_wire[95];
assign internal_wire[97] = ~internal_wire[96];
assign internal_wire[98] = ~internal_wire[97];
assign internal_wire[99] = ~internal_wire[98];
assign internal_wire[100] = ~internal_wire[99];
assign internal_wire[101] = ~internal_wire[100];
assign internal_wire[102] = ~internal_wire[101];
assign internal_wire[103] = ~internal_wire[102];
assign internal_wire[104] = ~internal_wire[103];
assign internal_wire[105] = ~internal_wire[104];
assign internal_wire[106] = ~internal_wire[105];
assign internal_wire[107] = ~internal_wire[106];
assign internal_wire[108] = ~internal_wire[107];
assign internal_wire[109] = ~internal_wire[108];
assign internal_wire[110] = ~internal_wire[109];
assign internal_wire[111] = ~internal_wire[110];
assign internal_wire[112] = ~internal_wire[111];
assign internal_wire[113] = ~internal_wire[112];
assign internal_wire[114] = ~internal_wire[113];
assign internal_wire[115] = ~internal_wire[114];
assign internal_wire[116] = ~internal_wire[115];
assign internal_wire[117] = ~internal_wire[116];
assign internal_wire[118] = ~internal_wire[117];
assign internal_wire[119] = ~internal_wire[118];
assign internal_wire[120] = ~internal_wire[119];
assign internal_wire[121] = ~internal_wire[120];
assign internal_wire[122] = ~internal_wire[121];
assign internal_wire[123] = ~internal_wire[122];
assign internal_wire[124] = ~internal_wire[123];
assign internal_wire[125] = ~internal_wire[124];
assign internal_wire[126] = ~internal_wire[125];
assign internal_wire[127] = ~internal_wire[126];
assign internal_wire[128] = ~internal_wire[127];
assign internal_wire[129] = ~internal_wire[128];
assign internal_wire[130] = ~internal_wire[129];
assign internal_wire[131] = ~internal_wire[130];
assign internal_wire[132] = ~internal_wire[131];
assign internal_wire[133] = ~internal_wire[132];
assign internal_wire[134] = ~internal_wire[133];
assign internal_wire[135] = ~internal_wire[134];
assign internal_wire[136] = ~internal_wire[135];
assign internal_wire[137] = ~internal_wire[136];
assign internal_wire[138] = ~internal_wire[137];
assign internal_wire[139] = ~internal_wire[138];
assign internal_wire[140] = ~internal_wire[139];
assign internal_wire[141] = ~internal_wire[140];
assign internal_wire[142] = ~internal_wire[141];
assign internal_wire[143] = ~internal_wire[142];
assign internal_wire[144] = ~internal_wire[143];
assign internal_wire[145] = ~internal_wire[144];
assign internal_wire[146] = ~internal_wire[145];
assign internal_wire[147] = ~internal_wire[146];
assign internal_wire[148] = ~internal_wire[147];
assign internal_wire[149] = ~internal_wire[148];
assign internal_wire[150] = ~internal_wire[149];
assign internal_wire[151] = ~internal_wire[150];
assign internal_wire[152] = ~internal_wire[151];
assign internal_wire[153] = ~internal_wire[152];
assign internal_wire[154] = ~internal_wire[153];
assign internal_wire[155] = ~internal_wire[154];
assign internal_wire[156] = ~internal_wire[155];
assign internal_wire[157] = ~internal_wire[156];
assign internal_wire[158] = ~internal_wire[157];

//should be an even number: the last internal_wire: 158 corresponds to 160 not gates
endmodule